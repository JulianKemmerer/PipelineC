-- See make_image_files.py
-- pipelinec_color : ../../../../pipelinec_color.jpg
(
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(15, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(13, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(13, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(13, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(13, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(15, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(12, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(13, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(13, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(13, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(9, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(13, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(14, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(14, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(13, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(13, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(13, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(13, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(11, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(12, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(15, 4), g => to_unsigned(14, 4), b => to_unsigned(13, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(15, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(15, 4), g => to_unsigned(14, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(12, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(11, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(0, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(2, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(2, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(1, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(2, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(2, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(1, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(0, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(0, 4), g => to_unsigned(4, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(4, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(5, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(4, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(1, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(3, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(2, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(6, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(15, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(13, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(4, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(3, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(3, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(3, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(5, 4), b => to_unsigned(1, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(7, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(14, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(4, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(4, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(2, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(11, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(4, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(4, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(10, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(10, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(10, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(12, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(13, 4), b => to_unsigned(12, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(12, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(13, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(10, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(13, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(11, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(13, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(5, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(3, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(5, 4), g => to_unsigned(5, 4), b => to_unsigned(4, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(11, 4), b => to_unsigned(11, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(10, 4), b => to_unsigned(10, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(10, 4), b => to_unsigned(9, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(8, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(12, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(9, 4), b => to_unsigned(7, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(11, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(10, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(8, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(9, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(8, 4), g => to_unsigned(8, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(7, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(7, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(5, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(5, 4)),
(r => to_unsigned(6, 4), g => to_unsigned(6, 4), b => to_unsigned(6, 4))
)
