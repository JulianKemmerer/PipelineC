-- See make_image_files.py
-- pipelinec_color : ../../../../pipelinec_color.jpg
(
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(15, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(13, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(13, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(13, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(13, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(15, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(12, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(13, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(13, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(13, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(9, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(13, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(14, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(14, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(13, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(13, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(13, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(13, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(11, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(12, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(15, 4), green => to_unsigned(14, 4), blue => to_unsigned(13, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(15, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(15, 4), green => to_unsigned(14, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(12, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(11, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(0, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(2, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(2, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(1, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(2, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(2, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(1, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(0, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(0, 4), green => to_unsigned(4, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(4, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(5, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(4, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(1, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(3, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(2, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(6, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(15, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(13, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(4, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(3, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(3, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(3, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(5, 4), blue => to_unsigned(1, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(7, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(14, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(4, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(4, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(2, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(11, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(4, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(4, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(10, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(10, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(10, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(12, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(13, 4), blue => to_unsigned(12, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(12, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(13, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(10, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(13, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(11, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(13, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(5, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(3, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(5, 4), green => to_unsigned(5, 4), blue => to_unsigned(4, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(11, 4), blue => to_unsigned(11, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(10, 4), blue => to_unsigned(10, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(10, 4), blue => to_unsigned(9, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(8, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(12, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(9, 4), blue => to_unsigned(7, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(11, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(10, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(8, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(9, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(8, 4), green => to_unsigned(8, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(7, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(7, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(5, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(5, 4)),
(red => to_unsigned(6, 4), green => to_unsigned(6, 4), blue => to_unsigned(6, 4))
)